-- iclk.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity iclk is
	port (
		iclk_clk       : out std_logic;        --    iclk.clk
		iclk_en_oscena : in  std_logic := '0'  -- iclk_en.oscena
	);
end entity iclk;

architecture rtl of iclk is
	component altera_int_osc is
		port (
			oscena : in  std_logic := 'X'; -- oscena
			clkout : out std_logic         -- clk
		);
	end component altera_int_osc;

begin

	int_osc_0 : component altera_int_osc
		port map (
			oscena => iclk_en_oscena, -- oscena.oscena
			clkout => iclk_clk        -- clkout.clk
		);

end architecture rtl; -- of iclk
