
module iclk (
	iclk_en_oscena,
	iclk_clk);	

	input		iclk_en_oscena;
	output		iclk_clk;
endmodule
